`ifndef _sixbitexp_incl
`define _sixbitexp_incl

module sixbitexp(ain, out, overflow);
    input[5:0] ain;
    output[5:0] out;
    output overflow;
    
endmodule

`endif